module omega(output [7:0]z, input [7:0]x);

assign
  z=x;
endmodule
